typedef enum logic [2:0] {OP_AND=3'h3, OP_ADD=3'h2, OP_XOR=3'h4, OP_MULT=3'h1, OP_NULL=3'h0} opcode;
`define OP_CODES
